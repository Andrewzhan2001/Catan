0
0 0 0 0 0 r h 12 B 19 B
0 0 0 0 0 r h 13 B 18 B
0 0 0 0 0 r h 14 B 17 B
0 0 0 0 0 r h 15 B 16 B
