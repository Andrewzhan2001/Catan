0
0 0 0 0 0 r h 12 B
0 0 0 0 0 r h 25 B
0 0 0 0 0 r h 21 B
0 0 0 0 0 r h 35 B 47 B
0 10 4 11 2 5 2 5 3 9 1 4 4 6 5 7 0 3 1 8 1 8 3 2 4 4 2 9 0 6 2 3 3 12 1 10 0 11
7
