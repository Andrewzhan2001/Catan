3
1 1 2 0 0 r h 24 B 3 B
1 0 0 0 0 r h 35 B 12 B
3 0 0 0 0 r h 19 B 36 B
0 0 3 1 1 r h 27 B 50 B
2 8 1 6 4 3 3 5 0 10 1 11 5 7 2 6 0 4 2 8 2 5 4 12 4 4 0 11 3 9 0 3 1 9 1 2 3 10
6
