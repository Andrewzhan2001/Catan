0
0 0 0 0 0 r h 10 B 1 B
0 0 1 0 1 r h 34 B 44 B
0 0 0 0 0 r h 7 B 20 B
0 0 0 0 1 r h 2 B 52 B
