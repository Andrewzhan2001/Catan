Blue
10 10 10 10 10 r h 24 B 1 B
10 10 10 10 11 r h 15 B 10 B
10 10 10 10 10 r h 3 B 50 B
10 10 10 10 10 r h 19 B 27 B
2 5 1 11 2 9 4 4 4 3 2 8 1 8 3 4 3 5 0 11 2 2 0 3 0 6 5 7 3 10 1 9 1 12 4 10 0 6
13
