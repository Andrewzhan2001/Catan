0
0 0 0 1 0 r h 1 B 8 B
0 0 0 2 0 r h 2 B 7 B
0 0 0 1 0 r h 3 B 6 B
0 0 0 0 0 r h 4 B 5 B
