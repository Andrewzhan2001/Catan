0
10 10 11 10 10 r h 33 B 12 B
10 10 10 10 10 r h 25 B 42 B
10 10 10 10 10 r h 3 B 41 B
10 11 10 10 10 r h 53 B 30 B
