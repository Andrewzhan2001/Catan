2
10 10 10 10 10 r h 12 B 33 B
10 11 10 10 10 r h 24 B 50 B
10 10 10 10 10 r h 35 B 2 B
10 10 10 10 10 r h 17 B 9 B
5 7 4 8 0 2 2 6 2 5 3 6 1 4 0 3 1 3 3 9 4 5 2 10 2 10 0 12 3 9 1 8 4 11 0 11 1 4
0
