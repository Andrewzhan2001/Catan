1
2 1 7 6 4 r 29 36 h 27 B 24 B
2 0 1 1 7 r 22 0 h 0 B 14 B
0 1 4 5 8 r h 40 B 38 B
0 1 4 5 8 r h 50 B 10 B
